module functionABC(
	input logic A,B,C,
	output logic F
);



and(F, A, B);

endmodule